module xor_gate(
    output c,
    input a,b
    );
    xor g1(c,a,b);
endmodule
