module xnor_gate(
    output c,
    input a,b
    );
    xnor g1(c,a,b);
endmodule
