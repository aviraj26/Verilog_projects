module nor_gate(
    output c,
    input a,b
    );
    nor g1(c,a,b);
endmodule
