module and_gate(
    output c,
    input a,b
    );
    and g1(c,a,b);
endmodule
