module or_gate(
    output c,
    input a,b
    );
    or g1(c,a,b);
endmodule
