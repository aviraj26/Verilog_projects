module nand_gate(
    output c,
    input a,b
    );
    nand g1(c,a,b);
endmodule
